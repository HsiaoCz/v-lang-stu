module main

fn main() {
	println("world")
}